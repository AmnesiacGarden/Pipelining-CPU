library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_signed.all;
use ieee.std_logic_unsigned.all;

--*****************************************************************************
--**** ENTITY BSHIFT8
--****
--**** Description: This design shifts 16-bit data 8 places either by logic
--****              shifts left or right, arithmetic shift right or rotate 
--****              right. It shifts only when the enable line is set high.
--****              Otherwise it passes the 16-bit data through unchanged
--**** Version    : 1.0
--**** Date       : 12/8/99
--**** Programmer : Jason Gorham
--*****************************************************************************
ENTITY bshift8 IS
    PORT(data                           : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
         enable                         : IN STD_LOGIC;
         operation                      : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
         result                         : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END ENTITY bshift8;

ARCHITECTURE shift8_behav OF bshift8 IS
BEGIN
    name : PROCESS(data, enable, operation) IS
    CONSTANT zero : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
    BEGIN
        IF(enable='1') THEN
            CASE operation IS
                -- shift left logic by 8
                WHEN "00" => 
                    result <= data(7 DOWNTO 0) & zero;

                --shift right logic by 8
                WHEN "01" =>
                    result <= zero & data(15 DOWNTO 8);
            
                --arithmetic shift right by 8
                WHEN "10" =>
                    IF(data(15)='1') THEN
                        result <= "11111111" & data(15 DOWNTO 8);
                    ELSE
                        result <= zero & data(15 DOWNTO 8);
                    END IF;
            
                --rotate right
                WHEN OTHERS =>
                    result <= data(7 DOWNTO 0) & data(15 DOWNTO 8);

            END CASE;   
        ELSE
            --Enable line is not set so let data pass through unchanged
            result <= data;
        END IF; 
    END PROCESS name;
END ARCHITECTURE shift8_behav;      

    
